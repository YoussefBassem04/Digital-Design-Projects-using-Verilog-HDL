module uart_tx(
    input clk, 
    input reset, 
    input [7:0] data_in, 
    input start, 
    output reg tx, 
    output reg busy
);

endmodule